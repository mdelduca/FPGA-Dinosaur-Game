
module keyboard(
	input wire clk,
	input wire PS2_clk,
	input wire PS2_data,
	input wire[10:0] data,
	input parity,
	input stop
	);
	



endmodule
